`define A_TO_B_WIDTH 8
`define B_TO_A_WIDTH 16
`define A_EXTRA_WIDTH 4
`define B_EXTRA_WIDTH 12
