`define A_EXTRA_WIDTH 4
`define B_EXTRA_WIDTH 12
`define A_TO_B_BITWIDTH 8 
`define B_TO_A_BITWIDTH 16

`define DATA_FROM_B_BITWIDTH `B_TO_A_BITWIDTH
`define DATA_TO_B_BITWIDTH   `A_TO_B_BITWIDTH
`define DATA_FROM_A_BITWIDTH `A_TO_B_BITWIDTH
`define DATA_TO_A_BITWIDTH   `B_TO_A_BITWIDTH
`define A_EXTRA_IN_BITWIDTH  `A_EXTRA_WIDTH
`define A_EXTRA_OUT_BITWIDTH `A_EXTRA_WIDTH
`define B_EXTRA_IN_BITWIDTH  `B_EXTRA_WIDTH
`define B_EXTRA_OUT_BITWIDTH `B_EXTRA_WIDTH
