// top -> module_a, module_b
`define A_TO_B_BITWIDTH 8 
`define B_TO_A_BITWIDTH 16

// module_a
`define DATA_FROM_B_BITWIDTH `B_TO_A_BITWIDTH
`define DATA_TO_B_BITWIDTH   `A_TO_B_BITWIDTH
`define A_EXTRA_IN_BITWIDTH  4
`define A_EXTRA_OUT_BITWIDTH 4

// module_b
`define B_EXTRA_IN_BITWIDTH  12
`define B_EXTRA_OUT_BITWIDTH 12
`define DATA_FROM_A_BITWIDTH `A_TO_B_BITWIDTH
`define DATA_TO_A_BITWIDTH   `B_TO_A_BITWIDTH